-- y'' + 